#This should contain the wrapper file
